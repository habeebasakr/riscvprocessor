module InstMem (input [5:0] addr , output [31:0] data_out);
 reg [7:0] mem [0:255];
 assign data_out ={mem[3+addr],mem[2+addr],mem[1+addr], mem[addr]};
 initial begin
//  {mem[3],mem[2],mem[1],mem[0]}=
{mem[3],mem[2],mem[1],mem[0]}     =32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0                          
{mem[7],mem[6],mem[5],mem[4]}  =32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0) x1=17                         
{mem[11],mem[10],mem[9],mem[8]}    =32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0) x2=9                          
{mem[15],mem[14],mem[13],mem[12]}  =32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0) x3=25                      
{mem[19],mem[18],mem[17],mem[16]}   =32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2 x4=25                  
{mem[23],mem[22],mem[21],mem[20]}   =32'b0_000000_00011_00100_000_0100_0_1100011 ; //beq x4, x3, L               
{mem[27],mem[26],mem[25],mem[24]}  =32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2                
{mem[31],mem[30],mem[29],mem[28]}  =32'b0000000_00010_00011_000_00101_0110011 ; //L: add x5,x3,x2 x5=34         
{mem[35],mem[34],mem[33],mem[32]}   =32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0) mem[3]=34        
{mem[39],mem[38],mem[37],mem[36]}   =32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0) x6=34            
{mem[43],mem[42],mem[41],mem[40]}   =32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1 x7=0           
{mem[47],mem[46],mem[45],mem[44]}   =32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2 x8=8           
{mem[51],mem[50],mem[49],mem[48]}   =32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2 x0=0           
{mem[55],mem[54],mem[53],mem[52]} =32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1 x9=17  
//{mem[59],mem[58],mem[57],mem[56]} 
//{mem[63],mem[62],mem[61],mem[60]}
//{mem[67],mem[66],mem[65],mem[64]} 
//{mem[71],mem[70],mem[69],mem[68]} 
//{mem[75],mem[74],mem[73],mem[72]}
//{mem[79],mem[78],mem[77],mem[76]}
//{mem[83],mem[82],mem[81],mem[80]}
//{mem[87],mem[86],mem[85],mem[84]}
//{mem[91],mem[90],mem[89],mem[88]}
//{mem[95],mem[94],mem[93],mem[92]}
//{mem[99],mem[98],mem[97],mem[96]}
//{mem[103],mem[102],mem[101],mem[100]}
//{mem[107],mem[106],mem[105],mem[104]}
//{mem[111],mem[110],mem[109],mem[108]}
//{mem[115],mem[114],mem[113],mem[112]}
//{mem[119],mem[118],mem[117],mem[116]}
end
endmodule 